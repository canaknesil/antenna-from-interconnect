-- MIT License

-- Copyright (c) 2022 Can Aknesil

-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:

-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.

-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.MATH_REAL.ALL;


entity transmitter_data_src is
    generic(rom_size: integer := 2048);
    Port ( addr : in STD_LOGIC_VECTOR (integer(ceil(log2(real(rom_size))))-1 downto 0);
           dout : out STD_LOGIC);
end transmitter_data_src;


architecture Behavioral of transmitter_data_src is

signal rom: std_logic_vector(rom_size-1 downto 0);

begin

-- Barker_13_13 followed by random bits, 4bit-BPSK (1000, 0010), length = 2048
--rom <= "10001000100010001000001000101000100000101000001010001000100010001000100000100010100010000010100000101000100010001000100010000010001010001000001010000010100010001000100010001000001000101000100000101000001010001000100010001000100000100010100010000010100000101000001000100010001000101000100000100010100000101000001000100010001000100010100010000010001010000010100000101000100010001000100000100010100010000010100000101000100010001000100010000010001010001000001010000010100000100010001000100010100010000010001010000010100000101000100010001000100000100010100010000010100000101000001000100010001000101000100000100010100000101000001010001000100010001000001000101000100000101000001010001000001000101000001000100010001010001000001010001000001010001000100010000010100010001000100010000010001000100010001010001000100010000010001000100010100010000010100010001000100000101000001010000010100010001000001000101000100010000010100000100010001010001000001010000010001010000010100010001000001000101000001000100010100000101000100000100010100000101000100000100010001000100010100010000010001010000010001010000010100000100010100010001000001000100010100010000010001010001000001010001000100000101000100010000010001010000010001010000010001000100010001010001000001010000010100010000010001000101000100000101000001000100010100010001000001000101000001000101000001010001000100000100010100000100010001010001000001000100010100010001000100000101000001000101000100000101000001010000010001000101000100000101000001010000010001010000010100010000010001000101000001000100010001000100010100000101000100010001000100000101000100010000010001010000010100010001000001000101000100000101000100000100010100010001000001000100010100010000010100010001000001000100010100000100010001010000010100000100010100000100010100010000010100000100010001000101000001010000010001000101000001000100010001010001000001000100010001010001000100010001000100010000010001000100010001010001000100000101000100000101000001000101000100000100010001010001000001010000010100010000010001010001000001010000010001000101000001010001000";

-- Barker_13_13 followed by random bits, 2bit-AM (10, 00), length = 2048
rom <= "10101010100000101000100010101010101000001010001000101010101010000010100010001010101010100000101000100010101010101000001010001000100000000000101000001000100000000000001010000010001000101010101000001010001000101010101010000010100010001000000000001010000010001000101010101000001010001000100000000000101000001000100010101010100000101000100010000010001010100010001000100010001000000000001000001000100000100010100000100000101010100000000000101000101010101000001010101010001010000010000010100010100000000010101000100010001000001010001000001010101010000000101010001000100000000000100000101000101000000010101010101000101010101000000010001000000000100010001000001000100000100000000000000010101000001010001000001000101000101000000000100000000010101000001010101010001010000010000010101010001010100000100000000000000010100010000010000010001000001010000010100000100010000000100000001000001010101010000010101010101010001010101000000000100000100000101010100010100000100010000010100010000010001000001010101010101010001000001000100010101000101010001010001000100010000000100010101010000000000000100010101010001010101010100010101000001010101010100000101000101010000010000010000000101000101010000000001000000000100010100010100000101000000010000010000000000010001000001000001010000000001000001000100010001010000000000000101000001000000010101000101010001010100010001000001010000000100010101010101010100000000010100010001010001000101010100010001010100000101010000010000000101010000010001010000000101000100000001000000000100000101000001000000000000010101000101000101010001010101010101010100010101000101010101000000000000010101000101010101010001000100010000010000000001000000000100010101000000010100000100010001000100010001010001000000000100000100010101000001010000010101000100010100000100000100000100000100000100010101000000000100000000000100000000010001010101010000000101010000000000000101010001000101000101010101010000000000010101010100000101000101010001000101010000000000000001000000010101000100000101010101000000000101000000000101010100000000010000010100000001000100000";

dout <= rom(conv_integer(addr));


end Behavioral;
